module adder_i140_o71 (a,b,r);
input [69:0] a,b;
output [70:0] r;

assign r = a+b;

endmodule
