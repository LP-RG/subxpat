module adder_i88_o45 (a,b,r);
input [43:0] a,b;
output [44:0] r;

assign r = a+b;

endmodule
