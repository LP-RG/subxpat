module adder_i172_o87 (a,b,r);
input [85:0] a,b;
output [86:0] r;

assign r = a+b;

endmodule
