module adder_i220_o111 (a,b,r);
input [109:0] a,b;
output [110:0] r;

assign r = a+b;

endmodule
