module adder_i188_o95 (a,b,r);
input [93:0] a,b;
output [94:0] r;

assign r = a+b;

endmodule
