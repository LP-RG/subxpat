module mul_i8_o8_lpp0_ppo1_et128_SOP1_pap50_iter1 (in0, in1, in2, in3, in4, in5, in6, in7, out0, out1, out2, out3, out4, out5, out6, out7);
//input/output declarations
input in0, in1, in2, in3, in4, in5, in6, in7;
output out0, out1, out2, out3, out4, out5, out6, out7;
//intact gates wires 
wire w_g106, w_g107, w_g108, w_g109, w_g110, w_g111, w_g112, w_g113, w_g114, w_g115, w_g116, w_g117, w_g118, w_g119, w_g120, w_g121, w_g122, w_g123, w_g124, w_g125, w_g126, w_g127, w_g128, w_g129, w_g130, w_g131, w_g132, w_g133, w_g134, w_g135, w_g136, w_g137, w_g138, w_g139, w_g140, w_g141, w_g142, w_g143, w_g144, w_g145, w_g146, w_g147, w_g148, w_g149, w_g150, w_g151, w_g152, w_g153, w_g154, w_g155, w_g156, w_g157, w_g158, w_g159, w_g160, w_g161, w_g162, w_g163, w_g164, w_g165, w_g166, w_g167, w_g168, w_g169, w_g170, w_g171, w_g172, w_g173, w_g174, w_g175, w_g176, w_g177, w_g178, w_g179, w_g180, w_g181, w_g182, w_g183, w_g184, w_g185, w_g186, w_g187, w_g188, w_g189, w_g190, w_g191, w_g192, w_g193, w_g194, w_g195, w_g196, w_g197, w_g198, w_g199, w_g200, w_g201, w_g202, w_g203, w_g204, w_g205, w_g206, w_g207, w_g208, w_g209, w_g210;
//annotated subgraph inputs
wire w_in7, w_in6, w_in5, w_in4, w_in3, w_in2, w_in1, w_in0;
//annotated subgraph outputs
wire w_g24, w_g28, w_g40, w_g44, w_g47, w_g66, w_g69, w_g73, w_g75, w_g87, w_g88, w_g92, w_g99, w_g101, w_g102, w_g103, w_g104, w_g105;
//json input wires
wire j_in0, j_in1, j_in2, j_in3, j_in4, j_in5, j_in6, j_in7;
//json model
wire p_o0_t0, p_o1_t0, p_o2_t0, p_o3_t0, p_o4_t0, p_o5_t0, p_o6_t0, p_o7_t0, p_o8_t0, p_o9_t0, p_o10_t0, p_o11_t0, p_o12_t0, p_o13_t0, p_o14_t0, p_o15_t0, p_o16_t0, p_o17_t0;
//subgraph inputs assigns
assign w_in7 = in7;
assign w_in6 = in6;
assign w_in5 = in5;
assign w_in4 = in4;
assign w_in3 = in3;
assign w_in2 = in2;
assign w_in1 = in1;
assign w_in0 = in0;
//mapping subgraph inputs to json inputs
assign j_in0 = w_in0;
assign j_in1 = w_in1;
assign j_in2 = w_in2;
assign j_in3 = w_in3;
assign j_in4 = w_in4;
assign j_in5 = w_in5;
assign j_in6 = w_in6;
assign j_in7 = w_in7;
//json model assigns (approximated/XPATed part)
assign p_o0_t0 = 1;
assign w_g24 = p_o0_t0;
assign p_o1_t0 = 1;
assign w_g28 = p_o1_t0;
assign w_g40 = 0;
assign w_g44 = 0;
assign w_g47 = 0;
assign w_g66 = 0;
assign w_g69 = 0;
assign w_g73 = 0;
assign w_g75 = 0;
assign p_o9_t0 = 1;
assign w_g87 = p_o9_t0;
assign p_o10_t0 = 1;
assign w_g88 = p_o10_t0;
assign p_o11_t0 = 1;
assign w_g92 = p_o11_t0;
assign p_o12_t0 = 1;
assign w_g99 = p_o12_t0;
assign w_g101 = 0;
assign w_g102 = 0;
assign w_g103 = 0;
assign p_o16_t0 = 1;
assign w_g104 = p_o16_t0;
assign p_o17_t0 = 1;
assign w_g105 = p_o17_t0;
// intact gates assigns
assign w_g106 = ~w_g101;
assign w_g107 = w_g75 & w_g102;
assign w_g108 = ~w_g102;
assign w_g109 = w_g103 & w_g66;
assign w_g110 = ~w_g103;
assign w_g111 = ~w_g104;
assign w_g112 = w_g105 & w_g99;
assign w_g113 = w_g106 & w_g104;
assign w_g114 = ~w_g107;
assign w_g115 = w_g108 & w_g69;
assign w_g116 = ~w_g109;
assign w_g117 = w_g110 & w_g73;
assign w_g118 = w_g111 & w_g101;
assign w_g119 = ~w_g112;
assign w_g120 = ~w_g113;
assign w_g121 = ~w_g115;
assign w_g122 = ~w_g117;
assign w_g123 = ~w_g118;
assign w_g124 = ~w_g119;
assign w_g125 = w_g121 & w_g114;
assign w_g126 = w_g116 & w_g122;
assign w_g127 = ~w_g122;
assign w_g128 = w_g123 & w_g120;
assign w_g129 = ~w_g125;
assign w_g130 = ~w_g126;
assign w_g131 = ~w_g128;
assign w_g132 = w_g129 & w_g24;
assign w_g133 = ~w_g129;
assign w_g134 = ~w_g130;
assign w_g135 = w_g131 & w_g28;
assign w_g136 = ~w_g131;
assign w_g137 = ~w_g132;
assign w_g138 = w_g133 & w_g40;
assign w_g139 = ~w_g135;
assign w_g140 = w_g136 & w_g44;
assign w_g141 = ~w_g138;
assign w_g142 = ~w_g140;
assign w_g143 = w_g137 & w_g141;
assign w_g144 = w_g141 & w_g114;
assign w_g145 = w_g139 & w_g142;
assign w_g146 = w_g142 & w_g120;
assign w_g147 = ~w_g143;
assign w_g148 = ~w_g144;
assign w_g149 = ~w_g145;
assign w_g150 = ~w_g146;
assign w_g151 = ~w_g147;
assign w_g152 = w_g92 & w_g148;
assign w_g153 = ~w_g148;
assign w_g154 = w_g149 & w_g122;
assign w_g155 = ~w_g149;
assign w_g156 = ~w_g150;
assign w_g157 = w_g151 & w_g150;
assign w_g158 = ~w_g152;
assign w_g159 = w_g153 & w_g88;
assign w_g160 = ~w_g154;
assign w_g161 = w_g127 & w_g155;
assign w_g162 = w_g156 & w_g147;
assign w_g163 = ~w_g157;
assign w_g164 = ~w_g159;
assign w_g165 = ~w_g161;
assign w_g166 = ~w_g162;
assign w_g167 = w_g163 & w_g158;
assign w_g168 = ~w_g163;
assign w_g169 = w_g164 & w_g158;
assign w_g170 = w_g160 & w_g165;
assign w_g171 = ~w_g165;
assign w_g172 = w_g166 & w_g163;
assign w_g173 = ~w_g167;
assign w_g174 = w_g168 & w_g164;
assign w_g175 = ~w_g169;
assign w_g176 = ~w_g170;
assign w_g177 = ~w_g172;
assign w_g178 = w_g173 & w_g164;
assign w_g179 = ~w_g174;
assign w_g180 = ~w_g175;
assign w_g181 = ~w_g176;
assign w_g182 = w_g177 & w_g165;
assign w_g183 = ~w_g177;
assign w_g184 = ~w_g178;
assign w_g185 = w_g179 & w_g158;
assign w_g186 = ~w_g182;
assign w_g187 = w_g183 & w_g171;
assign w_g188 = w_g184 & w_g119;
assign w_g189 = ~w_g185;
assign w_g190 = ~w_g187;
assign w_g191 = ~w_g188;
assign w_g192 = w_g124 & w_g189;
assign w_g193 = w_g190 & w_g163;
assign w_g194 = w_g186 & w_g190;
assign w_g195 = ~w_g192;
assign w_g196 = ~w_g193;
assign w_g197 = ~w_g194;
assign w_g198 = w_g191 & w_g195;
assign w_g199 = w_g195 & w_g99;
assign w_g200 = w_g196 & w_g175;
assign w_g201 = ~w_g196;
assign w_g202 = ~w_g197;
assign w_g203 = ~w_g198;
assign w_g204 = ~w_g199;
assign w_g205 = ~w_g200;
assign w_g206 = w_g180 & w_g201;
assign w_g207 = ~w_g203;
assign w_g208 = ~w_g206;
assign w_g209 = w_g205 & w_g208;
assign w_g210 = ~w_g209;
// output assigns
assign out0 = w_g47;
assign out1 = w_g87;
assign out2 = w_g134;
assign out3 = w_g181;
assign out4 = w_g202;
assign out5 = w_g210;
assign out6 = w_g207;
assign out7 = w_g204;
endmodule