module adder_i248_o125 (a,b,r);
input [123:0] a,b;
output [124:0] r;

assign r = a+b;

endmodule
