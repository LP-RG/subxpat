module adder_i156_o79 (a,b,r);
input [77:0] a,b;
output [78:0] r;

assign r = a+b;

endmodule
