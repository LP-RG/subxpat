module adder_i236_o119 (a,b,r);
input [117:0] a,b;
output [118:0] r;

assign r = a+b;

endmodule
