module adder_i124_o63 (a,b,r);
input [61:0] a,b;
output [62:0] r;

assign r = a+b;

endmodule
