module adder_i116_o59 (a,b,r);
input [57:0] a,b;
output [58:0] r;

assign r = a+b;

endmodule
