module adder_i244_o123 (a,b,r);
input [121:0] a,b;
output [122:0] r;

assign r = a+b;

endmodule
