module adder_i184_o93 (a,b,r);
input [91:0] a,b;
output [92:0] r;

assign r = a+b;

endmodule
