module adder_i176_o89 (a,b,r);
input [87:0] a,b;
output [88:0] r;

assign r = a+b;

endmodule
