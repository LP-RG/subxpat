module adder_i100_o51 (a,b,r);
input [49:0] a,b;
output [50:0] r;

assign r = a+b;

endmodule
