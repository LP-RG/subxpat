module adder_i72_o37 (a,b,r);
input [35:0] a,b;
output [36:0] r;

assign r = a+b;

endmodule
