module adder_i104_o53 (a,b,r);
input [51:0] a,b;
output [52:0] r;

assign r = a+b;

endmodule
