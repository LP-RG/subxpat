module adder_i192_o97 (a,b,r);
input [95:0] a,b;
output [96:0] r;

assign r = a+b;

endmodule
