module adder_i76_o39 (a,b,r);
input [37:0] a,b;
output [38:0] r;

assign r = a+b;

endmodule
