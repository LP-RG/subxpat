module adder_i168_o85 (a,b,r);
input [83:0] a,b;
output [84:0] r;

assign r = a+b;

endmodule
