module adder_i164_o83 (a,b,r);
input [81:0] a,b;
output [82:0] r;

assign r = a+b;

endmodule
