module adder_i200_o101 (a,b,r);
input [99:0] a,b;
output [100:0] r;

assign r = a+b;

endmodule
