module adder_i148_o75 (a,b,r);
input [73:0] a,b;
output [74:0] r;

assign r = a+b;

endmodule
