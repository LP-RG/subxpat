module adder_i196_o99 (a,b,r);
input [97:0] a,b;
output [98:0] r;

assign r = a+b;

endmodule
