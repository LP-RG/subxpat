module adder_i224_o113 (a,b,r);
input [111:0] a,b;
output [112:0] r;

assign r = a+b;

endmodule
