module adder_i112_o57 (a,b,r);
input [55:0] a,b;
output [56:0] r;

assign r = a+b;

endmodule
