module adder_i232_o117 (a,b,r);
input [115:0] a,b;
output [116:0] r;

assign r = a+b;

endmodule
