module adder_i160_o81 (a,b,r);
input [79:0] a,b;
output [80:0] r;

assign r = a+b;

endmodule
