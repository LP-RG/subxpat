module adder_i144_o73 (a,b,r);
input [71:0] a,b;
output [72:0] r;

assign r = a+b;

endmodule
