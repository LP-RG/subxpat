module adder_i84_o43 (a,b,r);
input [41:0] a,b;
output [42:0] r;

assign r = a+b;

endmodule
