module adder_i120_o61 (a,b,r);
input [59:0] a,b;
output [60:0] r;

assign r = a+b;

endmodule
