module adder_i92_o47 (a,b,r);
input [45:0] a,b;
output [46:0] r;

assign r = a+b;

endmodule
