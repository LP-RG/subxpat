module adder_i216_o109 (a,b,r);
input [107:0] a,b;
output [108:0] r;

assign r = a+b;

endmodule
