module adder_i132_o67 (a,b,r);
input [65:0] a,b;
output [66:0] r;

assign r = a+b;

endmodule
