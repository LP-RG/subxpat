module adder_i252_o127 (a,b,r);
input [125:0] a,b;
output [126:0] r;

assign r = a+b;

endmodule
