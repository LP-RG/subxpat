module adder_i212_o107 (a,b,r);
input [105:0] a,b;
output [106:0] r;

assign r = a+b;

endmodule
