module adder_i68_o35 (a,b,r);
input [33:0] a,b;
output [34:0] r;

assign r = a+b;

endmodule
