module adder_i108_o55 (a,b,r);
input [53:0] a,b;
output [54:0] r;

assign r = a+b;

endmodule
