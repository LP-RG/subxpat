module adder_i228_o115 (a,b,r);
input [113:0] a,b;
output [114:0] r;

assign r = a+b;

endmodule
