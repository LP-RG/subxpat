module adder_i240_o121 (a,b,r);
input [119:0] a,b;
output [120:0] r;

assign r = a+b;

endmodule
