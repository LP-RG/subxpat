module adder_i204_o103 (a,b,r);
input [101:0] a,b;
output [102:0] r;

assign r = a+b;

endmodule
