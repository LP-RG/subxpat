module adder_i208_o105 (a,b,r);
input [103:0] a,b;
output [104:0] r;

assign r = a+b;

endmodule
