module adder_i136_o69 (a,b,r);
input [67:0] a,b;
output [68:0] r;

assign r = a+b;

endmodule
