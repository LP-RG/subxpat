module adder_i80_o41 (a,b,r);
input [39:0] a,b;
output [40:0] r;

assign r = a+b;

endmodule
