module adder_i96_o49 (a,b,r);
input [47:0] a,b;
output [48:0] r;

assign r = a+b;

endmodule
