module adder_i152_o77 (a,b,r);
input [75:0] a,b;
output [76:0] r;

assign r = a+b;

endmodule
