module adder_i180_o91 (a,b,r);
input [89:0] a,b;
output [90:0] r;

assign r = a+b;

endmodule
