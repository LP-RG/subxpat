module adder_i256_o129 (a,b,r);
input [127:0] a,b;
output [128:0] r;

assign r = a+b;

endmodule
